// cat > counter.v << 'EOF'                                                                                                                                                      > module counter (                                                                                                                                                                                      >     input wire clk,                                                                                                                                                                                   >     input wire rst_n,                                                                                                                                                                                 >     input wire enable,                                                                                                                                                                                >     output reg [3:0] count,                                                                                                                                                                           >     output wire overflow                                                                                                                                                                              > );                                                                                                                                                                                                    >                                                                                                                                                                                                       > // Counter logic                                                                                                                                                                                      > always @(posedge clk or negedge rst_n) begin                                                                                                                                                          >     if (!rst_n) begin                                                                                                                                                                                 >         count <= 4'b0000;                                                                                                                                                                             >     end else if (enable) begin                                                                                                                                                                        >         count <= count + 1;                                                                                                                                                                           >     end                                                                                                                                                                                               > end                                                                                                                                                                                                   >                                                                                                                                                                                                       > // Overflow detection                                                                                                                                                                                 > assign overflow = (count == 4'b1111) & enable;                                                                                                                                                        >                                                                                                                                                                                                       > endmodule                                                                                                                                                                                             > EOF                     cat > counter.v << 'EOF'                                                                                                                                                      > module counter (                                                                                                                                                                                      >     input wire clk,                                                                                                                                                                                   >     input wire rst_n,                                                                                                                                                                                 >     input wire enable,                                                                                                                                                                                >     output reg [3:0] count,                                                                                                                                                                           >     output wire overflow                                                                                                                                                                              > );                                                                                                                                                                                                    >                                                                                                                                                                                                       > // Counter logic                                                                                                                                                                                      > always @(posedge clk or negedge rst_n) begin                                                                                                                                                          >     if (!rst_n) begin                                                                                                                                                                                 >         count <= 4'b0000;                                                                                                                                                                             >     end else if (enable) begin                                                                                                                                                                        >         count <= count + 1;                                                                                                                                                                           >     end                                                                                                                                                                                               > end                                                                                                                                                                                                   >                                                                                                                                                                                                       > // Overflow detection                                                                                                                                                                                 > assign overflow = (count == 4'b1111) & enable;                                                                                                                                                        >                                                                                                                                                                                                       > endmodule                                                 cat > counter.v << 'EOF'
module counter (
    input wire clk,
    input wire rst_n,
    input wire enable,
    output reg [3:0] count,
    output wire overflow
);

// Counter logic
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        count <= 4'b0000;
    end else if (enable) begin
        count <= count + 1;
    end
end

// Overflow detection
assign overflow = (count == 4'b1111) & enable;

endmodule
EOF                                                                                                                                         > EOF                     
